library verilog;
use verilog.vl_types.all;
entity pratica3 is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end pratica3;
